/usr/pack/umc-65-kgf/umc/ll/uk65lscllmvbbl/b03/lef/uk65lscllmvbbl.lef