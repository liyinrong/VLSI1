.SUBCKT MOMCAPS_SY_MMKF PLUS MINUS B
.ENDS

.SUBCKT MOMCAPS_AS_MMKF PLUS MINUS B
.ENDS

.SUBCKT MOMCAPS_SYMESH_MMKF PLUS1 MINUS1 PLUS2 MINUS2 B
.ENDS

.SUBCKT MOMCAPS_ASMESH_MMKF PLUS1 MINUS1 PLUS2 MINUS2 B
.ENDS

.SUBCKT MIMCAPS_20F_NWELL_RFKF PLUS MINUS NW PSUB
.ENDS

.SUBCKT MIMCAPS_20F_M1_RFKF PLUS MINUS PSUB
.ENDS

.SUBCKT MIMCAPS_20F_PSUB_RFKF PLUS MINUS PSUB
.ENDS

.SUBCKT VARDIOP_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT L_SLCR30K_RFVIL PLUS MINUS PSUB
.ENDS

.SUBCKT L_SQSK_RFVIL PLUS MINUS PSUB
.ENDS

.SUBCKT L_SY30K_RFVIL PLUS MINUS PSUB
.ENDS

.SUBCKT L_SYCT30K_RFVIL PLUS MINUS CT PSUB
.ENDS

.SUBCKT L_SLCR8K_RFVIL PLUS MINUS PSUB
.ENDS

.SUBCKT L_SY8K_RFVIL PLUS MINUS PSUB
.ENDS

.SUBCKT L_SYCT8K_RFVIL PLUS MINUS CT PSUB
.ENDS

.SUBCKT L_OCCTOUT_TRANS_RFVIL P1 P2 S1 S2 CTS PSUB
.ENDS

.SUBCKT L_SQ_TRANS_RFVIL P1 P2 S1 S2 PSUB
.ENDS

.SUBCKT L_SQCTIN_TRANS_RFVIL P1 P2 S1 S2 CTP PSUB
.ENDS

.SUBCKT L_SQCTOUT_TRANS_RFVIL P1 P2 S1 S2 CTS PSUB
.ENDS

.SUBCKT L_SQCTINOUT_TRANS_RFVIL P1 P2 S1 S2 CTP CTS PSUB
.ENDS

.SUBCKT MOMCAPS_Array_VP3_RFVCL PLUS MINUS NW PSUB
.ENDS

.SUBCKT MOMCAPS_Array_VP4_RFVCL PLUS MINUS NW PSUB
.ENDS

.SUBCKT MOMCAPS_Array_VP5_RFVCL PLUS MINUS SUB
.ENDS

.SUBCKT N_12_LLRVTRF D G S B
.ENDS

.SUBCKT N_12_LLHVTRF D G S B
.ENDS

.SUBCKT N_12_LLLVTRF D G S B
.ENDS

.SUBCKT N_18_LLRF D G S B
.ENDS

.SUBCKT N_25_LLRF D G S B
.ENDS

.SUBCKT N_33_LLRF D G S B
.ENDS

.SUBCKT N_BPW_12_LLRVTRF D G S B NW PSUB
.ENDS

.SUBCKT N_BPW_12_LLHVTRF D G S B NW PSUB
.ENDS

.SUBCKT N_BPW_12_LLLVTRF D G S B NW PSUB
.ENDS

.SUBCKT N_BPW_18_LLRF D G S B NW PSUB
.ENDS

.SUBCKT N_BPW_25_LLRF D G S B NW PSUB
.ENDS

.SUBCKT N_BPW_33_LLRF D G S B NW PSUB
.ENDS

.SUBCKT P_12_LLRVTRF D G S B PSUB
.ENDS

.SUBCKT P_12_LLHVTRF D G S B PSUB
.ENDS

.SUBCKT P_12_LLLVTRF D G S B PSUB
.ENDS

.SUBCKT P_18_LLRF D G S B PSUB
.ENDS

.SUBCKT P_25_LLRF D G S B PSUB
.ENDS

.SUBCKT P_33_LLRF D G S B PSUB
.ENDS

.SUBCKT RNHR_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT RNHR_NW_LLRF PLUS MINUS NW PSUB
.ENDS

.SUBCKT RNNPO_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT RNNPO_NW_LLRF PLUS MINUS NW PSUB
.ENDS

.SUBCKT RNPPO_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT RNPPO_NW_LLRF PLUS MINUS NW PSUB
.ENDS

.SUBCKT VARMIS_12_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT VARMIS_18_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT VARMIS_25_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT VARMIS_33_LLRF PLUS MINUS PSUB
.ENDS

.SUBCKT PAD_RF PLUS PSUB
.ENDS
