/usr/pack/umc-65-kgf/dz/encounter/13/u65ll_8m1t0f1u.lef