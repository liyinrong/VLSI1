/usr/pack/umc-65-kgf/umc/ll/u065gioll25mvir/b04/lef.dz/u065gioll25mvir_8m1t0f1u.lef